module wb_stage( input  wire [31:0] new_register_data,
                    input  wire is_write,
                    input  wire [3:0]  data_register_d);


endmodule
